`ifndef ADDER_TYPES
`define ADDER_TYPES

`endif